


entity contring00 is
	port(
		clkcr: in std_logic;
		ecr: in std_logic
		outcr: out std_logic_vector(3 downto 0)
	);
	
end contring00;